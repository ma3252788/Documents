library verilog;
use verilog.vl_types.all;
entity test_7180_v is
end test_7180_v;
