`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:11:10 03/17/2017 
// Design Name: 
// Module Name:    I2C_CTRL7179 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module I2C_CTRL7179(clk,rst,din,ack,err,rty,sel,
							cyc,stb,we,dout,adr,Finish
    );
	 
	
	input clk;
	input rst;
	input [7:0] din;
	input ack,

endmodule
