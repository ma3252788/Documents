library verilog;
use verilog.vl_types.all;
entity tst_dpram_v is
end tst_dpram_v;
